module new_module();

endmodule

